// sigmoid activation using fixed-point LUT approximation
module activation_sigmoid #(
    parameter WIDTH = 32,
    parameter FRAC_BITS = 16,
    parameter LUT_SIZE = 256
)(
    input  logic signed [WIDTH-1:0] in_data,
    output logic [WIDTH-1:0]         out_data
);

    logic [WIDTH-1:0] sigmoid_lut [0:LUT_SIZE-1];

    logic [7:0] lut_index;
    always_comb begin
        if (in_data < -((WIDTH>(FRAC_BITS+7)) ? (1 << (FRAC_BITS + 7)) : (1 << (WIDTH-1)))) 
            lut_index = 0;
        else if (in_data > ((WIDTH>(FRAC_BITS+7)) ? (1 << (FRAC_BITS + 7)) : (1 << (WIDTH-1))))
            lut_index = LUT_SIZE-1;
        else
            lut_index = (in_data >>> (FRAC_BITS - 8)) + (LUT_SIZE / 2); // Center LUT at 0
    end

    // lut output
    assign out_data = sigmoid_lut[lut_index];

    // initialise lut
    initial begin
        sigmoid_lut[0] = 22;
        sigmoid_lut[1] = 23;
        sigmoid_lut[2] = 25;
        sigmoid_lut[3] = 27;
        sigmoid_lut[4] = 28;
        sigmoid_lut[5] = 30;
        sigmoid_lut[6] = 32;
        sigmoid_lut[7] = 34;
        sigmoid_lut[8] = 36;
        sigmoid_lut[9] = 39;
        sigmoid_lut[10] = 41;
        sigmoid_lut[11] = 44;
        sigmoid_lut[12] = 47;
        sigmoid_lut[13] = 50;
        sigmoid_lut[14] = 53;
        sigmoid_lut[15] = 56;
        sigmoid_lut[16] = 60;
        sigmoid_lut[17] = 64;
        sigmoid_lut[18] = 68;
        sigmoid_lut[19] = 72;
        sigmoid_lut[20] = 77;
        sigmoid_lut[21] = 82;
        sigmoid_lut[22] = 87;
        sigmoid_lut[23] = 93;
        sigmoid_lut[24] = 99;
        sigmoid_lut[25] = 105;
        sigmoid_lut[26] = 112;
        sigmoid_lut[27] = 119;
        sigmoid_lut[28] = 127;
        sigmoid_lut[29] = 135;
        sigmoid_lut[30] = 144;
        sigmoid_lut[31] = 153;
        sigmoid_lut[32] = 163;
        sigmoid_lut[33] = 174;
        sigmoid_lut[34] = 185;
        sigmoid_lut[35] = 197;
        sigmoid_lut[36] = 210;
        sigmoid_lut[37] = 223;
        sigmoid_lut[38] = 238;
        sigmoid_lut[39] = 253;
        sigmoid_lut[40] = 269;
        sigmoid_lut[41] = 287;
        sigmoid_lut[42] = 305;
        sigmoid_lut[43] = 325;
        sigmoid_lut[44] = 346;
        sigmoid_lut[45] = 368;
        sigmoid_lut[46] = 392;
        sigmoid_lut[47] = 417;
        sigmoid_lut[48] = 444;
        sigmoid_lut[49] = 472;
        sigmoid_lut[50] = 503;
        sigmoid_lut[51] = 535;
        sigmoid_lut[52] = 569;
        sigmoid_lut[53] = 606;
        sigmoid_lut[54] = 645;
        sigmoid_lut[55] = 686;
        sigmoid_lut[56] = 730;
        sigmoid_lut[57] = 777;
        sigmoid_lut[58] = 826;
        sigmoid_lut[59] = 879;
        sigmoid_lut[60] = 935;
        sigmoid_lut[61] = 995;
        sigmoid_lut[62] = 1058;
        sigmoid_lut[63] = 1125;
        sigmoid_lut[64] = 1197;
        sigmoid_lut[65] = 1273;
        sigmoid_lut[66] = 1354;
        sigmoid_lut[67] = 1440;
        sigmoid_lut[68] = 1531;
        sigmoid_lut[69] = 1627;
        sigmoid_lut[70] = 1730;
        sigmoid_lut[71] = 1839;
        sigmoid_lut[72] = 1954;
        sigmoid_lut[73] = 2077;
        sigmoid_lut[74] = 2207;
        sigmoid_lut[75] = 2344;
        sigmoid_lut[76] = 2491;
        sigmoid_lut[77] = 2645;
        sigmoid_lut[78] = 2809;
        sigmoid_lut[79] = 2983;
        sigmoid_lut[80] = 3167;
        sigmoid_lut[81] = 3361;
        sigmoid_lut[82] = 3567;
        sigmoid_lut[83] = 3785;
        sigmoid_lut[84] = 4015;
        sigmoid_lut[85] = 4258;
        sigmoid_lut[86] = 4515;
        sigmoid_lut[87] = 4786;
        sigmoid_lut[88] = 5071;
        sigmoid_lut[89] = 5373;
        sigmoid_lut[90] = 5691;
        sigmoid_lut[91] = 6025;
        sigmoid_lut[92] = 6377;
        sigmoid_lut[93] = 6748;
        sigmoid_lut[94] = 7137;
        sigmoid_lut[95] = 7546;
        sigmoid_lut[96] = 7975;
        sigmoid_lut[97] = 8425;
        sigmoid_lut[98] = 8897;
        sigmoid_lut[99] = 9391;
        sigmoid_lut[100] = 9907;
        sigmoid_lut[101] = 10446;
        sigmoid_lut[102] = 11009;
        sigmoid_lut[103] = 11596;
        sigmoid_lut[104] = 12207;
        sigmoid_lut[105] = 12842;
        sigmoid_lut[106] = 13502;
        sigmoid_lut[107] = 14187;
        sigmoid_lut[108] = 14897;
        sigmoid_lut[109] = 15632;
        sigmoid_lut[110] = 16391;
        sigmoid_lut[111] = 17174;
        sigmoid_lut[112] = 17981;
        sigmoid_lut[113] = 18811;
        sigmoid_lut[114] = 19664;
        sigmoid_lut[115] = 20538;
        sigmoid_lut[116] = 21433;
        sigmoid_lut[117] = 22348;
        sigmoid_lut[118] = 23281;
        sigmoid_lut[119] = 24231;
        sigmoid_lut[120] = 25197;
        sigmoid_lut[121] = 26177;
        sigmoid_lut[122] = 27169;
        sigmoid_lut[123] = 28172;
        sigmoid_lut[124] = 29184;
        sigmoid_lut[125] = 30203;
        sigmoid_lut[126] = 31227;
        sigmoid_lut[127] = 32254;
        sigmoid_lut[128] = 33282;
        sigmoid_lut[129] = 34309;
        sigmoid_lut[130] = 35333;
        sigmoid_lut[131] = 36352;
        sigmoid_lut[132] = 37364;
        sigmoid_lut[133] = 38367;
        sigmoid_lut[134] = 39359;
        sigmoid_lut[135] = 40339;
        sigmoid_lut[136] = 41305;
        sigmoid_lut[137] = 42255;
        sigmoid_lut[138] = 43188;
        sigmoid_lut[139] = 44103;
        sigmoid_lut[140] = 44998;
        sigmoid_lut[141] = 45872;
        sigmoid_lut[142] = 46725;
        sigmoid_lut[143] = 47555;
        sigmoid_lut[144] = 48362;
        sigmoid_lut[145] = 49145;
        sigmoid_lut[146] = 49904;
        sigmoid_lut[147] = 50639;
        sigmoid_lut[148] = 51349;
        sigmoid_lut[149] = 52034;
        sigmoid_lut[150] = 52694;
        sigmoid_lut[151] = 53329;
        sigmoid_lut[152] = 53940;
        sigmoid_lut[153] = 54527;
        sigmoid_lut[154] = 55090;
        sigmoid_lut[155] = 55629;
        sigmoid_lut[156] = 56145;
        sigmoid_lut[157] = 56639;
        sigmoid_lut[158] = 57111;
        sigmoid_lut[159] = 57561;
        sigmoid_lut[160] = 57990;
        sigmoid_lut[161] = 58399;
        sigmoid_lut[162] = 58788;
        sigmoid_lut[163] = 59159;
        sigmoid_lut[164] = 59511;
        sigmoid_lut[165] = 59845;
        sigmoid_lut[166] = 60163;
        sigmoid_lut[167] = 60465;
        sigmoid_lut[168] = 60750;
        sigmoid_lut[169] = 61021;
        sigmoid_lut[170] = 61278;
        sigmoid_lut[171] = 61521;
        sigmoid_lut[172] = 61751;
        sigmoid_lut[173] = 61969;
        sigmoid_lut[174] = 62175;
        sigmoid_lut[175] = 62369;
        sigmoid_lut[176] = 62553;
        sigmoid_lut[177] = 62727;
        sigmoid_lut[178] = 62891;
        sigmoid_lut[179] = 63045;
        sigmoid_lut[180] = 63192;
        sigmoid_lut[181] = 63329;
        sigmoid_lut[182] = 63459;
        sigmoid_lut[183] = 63582;
        sigmoid_lut[184] = 63697;
        sigmoid_lut[185] = 63806;
        sigmoid_lut[186] = 63909;
        sigmoid_lut[187] = 64005;
        sigmoid_lut[188] = 64096;
        sigmoid_lut[189] = 64182;
        sigmoid_lut[190] = 64263;
        sigmoid_lut[191] = 64339;
        sigmoid_lut[192] = 64411;
        sigmoid_lut[193] = 64478;
        sigmoid_lut[194] = 64541;
        sigmoid_lut[195] = 64601;
        sigmoid_lut[196] = 64657;
        sigmoid_lut[197] = 64710;
        sigmoid_lut[198] = 64759;
        sigmoid_lut[199] = 64806;
        sigmoid_lut[200] = 64850;
        sigmoid_lut[201] = 64891;
        sigmoid_lut[202] = 64930;
        sigmoid_lut[203] = 64967;
        sigmoid_lut[204] = 65001;
        sigmoid_lut[205] = 65033;
        sigmoid_lut[206] = 65064;
        sigmoid_lut[207] = 65092;
        sigmoid_lut[208] = 65119;
        sigmoid_lut[209] = 65144;
        sigmoid_lut[210] = 65168;
        sigmoid_lut[211] = 65190;
        sigmoid_lut[212] = 65211;
        sigmoid_lut[213] = 65231;
        sigmoid_lut[214] = 65249;
        sigmoid_lut[215] = 65267;
        sigmoid_lut[216] = 65283;
        sigmoid_lut[217] = 65298;
        sigmoid_lut[218] = 65313;
        sigmoid_lut[219] = 65326;
        sigmoid_lut[220] = 65339;
        sigmoid_lut[221] = 65351;
        sigmoid_lut[222] = 65362;
        sigmoid_lut[223] = 65373;
        sigmoid_lut[224] = 65383;
        sigmoid_lut[225] = 65392;
        sigmoid_lut[226] = 65401;
        sigmoid_lut[227] = 65409;
        sigmoid_lut[228] = 65417;
        sigmoid_lut[229] = 65424;
        sigmoid_lut[230] = 65431;
        sigmoid_lut[231] = 65437;
        sigmoid_lut[232] = 65443;
        sigmoid_lut[233] = 65449;
        sigmoid_lut[234] = 65454;
        sigmoid_lut[235] = 65459;
        sigmoid_lut[236] = 65464;
        sigmoid_lut[237] = 65468;
        sigmoid_lut[238] = 65472;
        sigmoid_lut[239] = 65476;
        sigmoid_lut[240] = 65480;
        sigmoid_lut[241] = 65483;
        sigmoid_lut[242] = 65486;
        sigmoid_lut[243] = 65489;
        sigmoid_lut[244] = 65492;
        sigmoid_lut[245] = 65495;
        sigmoid_lut[246] = 65497;
        sigmoid_lut[247] = 65500;
        sigmoid_lut[248] = 65502;
        sigmoid_lut[249] = 65504;
        sigmoid_lut[250] = 65506;
        sigmoid_lut[251] = 65508;
        sigmoid_lut[252] = 65509;
        sigmoid_lut[253] = 65511;
        sigmoid_lut[254] = 65513;
        sigmoid_lut[255] = 65514;
    end

endmodule
