module multiplier #(parameter WIDTH = 32) (
    input logic [WIDTH-1:0] a,
    input logic [WIDTH-1:0] b,
    output logic [WIDTH-1:0] product
);

    assign product = a * b;

endmodule
